--Engineer      : Yinghao Li
--Created       : 11/19/2018
--Last Modified : 11/19/2018
--Name of file  : encoder_pkg.vhd
--Description   : Implementation of convolutional encoder

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

package encoder_pkg is

  constant STATE_NUM : integer := 10; -- TODO: subject to change

end encoder_pkg;

